module ALU
(   
    input  wire        clk,
    input  wire        rst,
    input  wire [31:0] a_in,
    input  wire [31:0] b_in,
    input  wire [3:0]  alu_control_in,
    input  wire        tick_idex,
    input  wire [31:0] pc,
    output reg  [31:0] alu_result,
    output reg         zero,
    output reg         cout,
    output reg         overflow
);




reg [32:0] result_temp;
reg [31:0] a;
reg [31:0] b;
reg [3:0]  alu_control;
reg [31:0] pc_reg;

always @(posedge clk) begin
    if(rst) begin
        result_temp = 33'd0;
        alu_result = 32'd0;
        zero = 1'b1;
        cout = 1'b0;
        overflow = 1'b0;
        a <= 32'd0;
        b <= 32'd0;
        alu_control <= 4'd0;
        pc_reg <= 32'd0;
    end
    else if(tick_idex) begin
        a <= a_in;
        b <= b_in;
        alu_control <= alu_control_in;
        pc_reg <= pc;
        result_temp <= 33'd0;
        alu_result <= 32'd0;
        zero <= 1'b1;
        cout <= 1'b0;
        overflow <= 1'b0;
    end
    else begin
        case (alu_control)
            4'b0000: begin   // ADD
                result_temp <= a + b;
                zero <= (result_temp == 33'd0);
                cout <= result_temp[32];
                overflow <= ((a[31] == b[31]) && (result_temp[31] != a[31]));
                alu_result <= result_temp[31:0];
            end
            4'b0001: begin   // SUB
                result_temp <= a + {1'b0, ~b} + 33'b1;
                zero <= (result_temp == 33'd0);
                cout <= result_temp[32];
                overflow <= ((a[31] != b[31]) && (result_temp[31] != a[31]));
                alu_result <= result_temp[31:0];
            end
            4'b0010: begin // Not A
                result_temp <= {1'b0, ~a};
                zero <= (result_temp == 33'd0);
                cout <= result_temp[32];
                overflow <= 1'b0;
                alu_result <= result_temp[31:0];
            end
            4'b0011: begin // A AND B
                result_temp <= {1'b0, a & b};
                zero <= (result_temp == 33'd0);
                cout <= result_temp[32];
                overflow <= 1'b0;
                alu_result <= result_temp[31:0];
            end
            4'b0100: begin // A OR B
                result_temp <= {1'b0, a | b};
                zero <= (result_temp == 33'd0);
                cout <= result_temp[32];
                overflow <= 1'b0;
                alu_result <= result_temp[31:0];
            end
            4'b0101: begin // A XOR B
                result_temp <= {1'b0, a ^ b};
                zero <= (result_temp == 33'd0);
                cout <= result_temp[32];
                overflow <= 1'b0;
                alu_result <= result_temp[31:0];
            end
            4'b0110: begin // SLT
                result_temp <= a + ({1'b0, ~b} + 33'b1);
                zero <= (result_temp == 33'd0);
                cout <= result_temp[32];
                overflow <= ((a[31] != b[31]) && (result_temp[31] != a[31]));
                alu_result <= ((((a[31] != b[31]) && (result_temp[31] != a[31])) ? ~result_temp[31] : result_temp[31]) && (result_temp[31] != 1'b0)) ? 32'd1 : 32'd0;
            end
            4'b0111: begin // EQU
                result_temp <= a + ({1'b0, ~b} + 33'b1);
                zero <= (result_temp == 33'd0);
                cout <= result_temp[32];
                overflow <= 1'b0;
                alu_result <= {result_temp == 33'd0 ? 32'd1 : 32'd0};
            end
            4'b1000: begin // SLL
                result_temp <= a << b[4:0];
                zero <= (result_temp == 33'd0);
                cout <= result_temp[32];
                overflow <= 1'b0;
                alu_result <= result_temp[31:0];
            end
            4'b1001: begin // SLTU
                result_temp <= a + ({1'b0, ~b} + 33'b1);
                zero <= (result_temp == 33'd0);
                cout <= result_temp[32];
                overflow <= ((a[31] != b[31]) && (result_temp[31] != a[31]));
                alu_result <= result_temp[31] && a[31] == 0 ? 32'd1 : 32'd0;
            end
            4'b1010: begin // SRL
                result_temp <= a >> b[4:0];
                zero <= (result_temp == 33'd0);
                cout <= result_temp[32];
                overflow <= 1'b0;
                alu_result <= result_temp[31:0];
            end
            4'b1011: begin // SRA
                result_temp <= ($signed(a)) >>> b[4:0];
                zero <= (result_temp == 33'd0);
                cout <= result_temp[32];
                overflow <= 1'b0;
                alu_result <= result_temp[31:0];
            end
            4'b1100: begin // LUI
                result_temp <= b ;
                zero <= (result_temp == 33'd0);
                cout <= result_temp[32];
                overflow <= 1'b0;
                alu_result <= result_temp[31:0];
            end
            4'b1101: begin // AUIPC
                result_temp <= pc_reg + b;
                zero <= (result_temp == 33'd0);
                cout <= result_temp[32];
                overflow <= 1'b0;
                alu_result <= result_temp[31:0];
            end
            default: begin
                result_temp <= 33'd0;
                alu_result <= 32'd0;
                zero <= 1'b1;
                cout <= 1'b0;
                overflow <= 1'b0;
            end
        endcase
    end
end





endmodule


