module Opcode_ctrl (
    input  wire [6:0] funct7,
    output wire       branch,
    output wire       mem_read,
    output wire       mem2reg,
    output wire       alop,
    output wire       mem_write,
    output wire       alu_src,
    output wire       reg_write
);






endmodule