module top (
    input  wire        clk,
    input  wire        rst,
    input  wire        pc_write
);

    // Instantiate your CPU components here
    // For example, ALU, Register File, Control Unit, etc.

endmodule